import uvm_pkg::*;
`include "uvm_macros.svh"

`include "interface.sv"
`include "transaction.sv"
`include "sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"
